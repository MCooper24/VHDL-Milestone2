--------- Students: Martin Cooper & Antonio Tembo ------
-------------- Numbers: UP736129 & UP504815 ------------
---------------- Module: THIRD - Channel 0 -------------

library ieee;																			
use ieee.std_logic_1164.all;				
use ieee.numeric_std.all;	

entity T17_M2_ChannelZero is
end T17_M2_ChannelZero;

architecture Behavioral of T17_M2_ChannelZero is

begin

end Behavioral;