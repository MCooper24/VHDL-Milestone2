--------- Students: Martin Cooper & Antonio Tembo ------
-------------- Numbers: UP736129 & UP504815 ------------
---------------- Module: FOURTH - Channel 1 ------------

library ieee;																			
use ieee.std_logic_1164.all;				
use ieee.numeric_std.all;	

entity T17_M2_ChannelOne is
end T17_M2_ChannelOne;

architecture Behavioral of T17_M2_ChannelOne is

begin

end Behavioral;